//-----------------------------------------------------------------
//--------------------------------------------------------------------
// Small RISC-V
// ALU, DATAPATH, CONTROL UNIT, IF/ID, ID/EX, EX/MEM, MEM/WB, NO STALL UNIT
//--------------------------------------------------------------------

module RISCV_CLOCK(clock);
    // OP-CODES
    parameter BEQ = 7'
