`include "DEFS.sv"

module adder #(
  parameter WIDTH = 32) //delay
  (
    input  [WIDTH-1:0] in1,
    input  [WIDTH-1:0] in2,
    output [WIDTH-1:0] result
);



endmodule
